library ieee;

use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.VIDEO_CONSTANTS.all;
use work.My_component_pkg.all;
---------------------------------------------------------------
-- ?????? ?????????? ?????????????
-- ???????? ?????? ? 3 ????????? ???????????? ??? / LVDS (1-2-4 ?????) / CSI (1 ?????)
-- ? ??????????? ?? mode_IMAGE_SENSOR (use work.VIDEO_CONSTANTS.all ) ????? ???????? ????? ?????????
-- mode_IMAGE_SENSOR (3 downto 0) = 0 CSI - 1 ?????
-- mode_IMAGE_SENSOR (3 downto 0) = 1 LVDS - 1 ?????
-- mode_IMAGE_SENSOR (3 downto 0) = 2 LVDS - 2 ?????
-- mode_IMAGE_SENSOR (3 downto 0) = 3 LVDS - 4 ?????
-- ??????????? ?????? ???????????? bit_data_imx 12 / 10 / 8 bit

-- mode_IMAGE_SENSOR (7 downto 4) = 0 B/W
-- mode_IMAGE_SENSOR (7 downto 4) = 1 COLOR

-- mode_generator ?????????? ??? ?????? ??? ????????
-- ??????? 4 ???? ??????? ?? ??? ???????, ??????? ?? ????????????
-- 	[7..4]						[3..0]
-- 	????? ????????				0 ???????????? ???? ?? ???????????
-- 	????? ????????				1 ???????????? ???? ?? ?????????
-- 	none							2 ???????????? ?????? ?? ?????? ???????? SMPTE
-- 	?????? ??????				3 ????????? ????
-- 	????????????? ?????		4 ??????? ?????? (color bar)
-- 	none							5 ?????? ?? ?????
--------------------------------------------------------------
--------------------------------------------------------------
-- ?????? PLL ??? ????????? ?????????????
-- ??? 2200?1250 50p ?????????? ??????? (PixFreq)  137.5 ???
-- ??? 2200?1125 30p ?????????? ??????? (PixFreq)  74.25 ???
-- ??? ?????????? ??????? > 74.25 ??? ?????? ??????????? CSI-2/ LVDS ?? 1 ?????
--       mode                        SerFreq
-- CSI      8 bit       PixFreq*4      = 297 ???
-- LVDS_1ch 8 bit       PixFreq*4      = 297 ???
-- LVDS_1ch 10 bit      PixFreq*5      = 371.25 ???
-- LVDS_1ch 12 bit      PixFreq*6      = 445.5 ???
-- LVDS_2ch 8 bit       PixFreq*4 /2   = 148.5 ???
-- LVDS_2ch 10 bit      PixFreq*5 /2   = 185.625 ???
-- LVDS_2ch 12 bit      PixFreq*6 /2   = 222.75 ???
-- LVDS_4ch 8 bit       PixFreq*4 /4   = 74.25 ???
-- LVDS_4ch 10 bit      PixFreq*5 /4   = 92.8125 ???
-- LVDS_4ch 12 bit      PixFreq*6 /4   = 111.375 ???
--------------------------------------------------------------

entity IMAGE_SENSOR_SIM_new is
port (
		--??????? ???????--	
	CLK					: in std_logic;  												-- ???????? 
	mode_generator		: in std_logic_vector (7 downto 0);						-- ??????? ??????????
		--???????? ???????--	
	XVS_Imx_Sim			: out std_logic; 												-- ?????????????
	XHS_Imx_Sim			: out std_logic; 												-- ?????????????
	DATA_IS_PAR			: out	std_logic_vector (bit_data_imx-1 downto 0);	-- ???????? ??????
	DATA_IS_LVDS_ch_n	: out	std_logic_vector (3 downto 0);					-- ???????? ?????? ? ?????? 1
	DATA_IS_CSI			: out	std_logic; 												-- ???????? ?????? CSI
	CLK_DDR				: out std_logic		
		);
end IMAGE_SENSOR_SIM_new;

architecture beh of IMAGE_SENSOR_SIM_new is 

----------------------------------------------------------------------
-- PLL_SIM_IS entity declaration
----------------------------------------------------------------------
component PLL_SIM_IS is
port( POWERDOWN : in    std_logic;
		CLKA      : in    std_logic;
		LOCK      : out   std_logic;
		GLA       : out   std_logic
		);
end component;
----------------------------------------------------------------------
-- PLL_SIM_IS entity declaration
----------------------------------------------------------------------
component PLL_SIM_IS_1 is
port( POWERDOWN : in    std_logic;
		CLKA      : in    std_logic;
		LOCK      : out   std_logic;
		GLA       : out   std_logic;
		GLB       : out   std_logic;
		GLC       : out   std_logic
		);
end component;

signal PLL_POWERDOWN_N	: std_logic;			
signal CLK_IS_pix			: std_logic;			
signal CLK_IS_DDR_0		: std_logic;			
signal CLK_IS_DDR_1		: std_logic;			
signal CLK_IS_DDR_2		: std_logic;			
signal locked_pll_0		: std_logic;
signal locked_pll_1		: std_logic;
signal main_enable		: std_logic;
signal main_reset			: std_logic;
signal locked_pll_q		: std_logic_vector(31 downto 0);
	
----------------------------------------------------------------------

----------------------------------------------------------------------
-- ?????? ????????? ???????????? ?? ????????????? ? ???????????? ????
----------------------------------------------------------------------
component IS_SIM_Paralell is
generic  (
	PixPerLine_is			: integer;
	HsyncShift_is			: integer;
	ActivePixPerLine_is	: integer;
	HsyncWidth_is			: integer;
	LinePerFrame_is		: integer;
	VsyncShift_is			: integer;
	ActiveLine_is			: integer;
	VsyncWidth_is			: integer
);
port (
		--??????? ???????--	
	CLK					: in std_logic;  												-- ???????? 
	main_reset			: in std_logic;  												-- main_reset
	main_enable			: in std_logic;  												-- main_enable
	mode_generator		: in std_logic_vector (7 downto 0);						--??????? ??????
		--???????? ???????--	
	qout_V_out			: out std_logic_vector (bit_strok-1 downto 0);		-- 
	qout_clk_out		: out std_logic_vector (bit_pix-1 downto 0 );		-- 
	XVS_Imx_Sim			: out std_logic; 												-- ?????????????
	XHS_Imx_Sim			: out std_logic; 												-- ?????????????
	DATA_IS_pix_ch_1	: out  std_logic_vector (bit_data_imx-1 downto 0);	-- ???????? ??????
	DATA_IS_pix_ch_2	: out  std_logic_vector (bit_data_imx-1 downto 0);	-- ???????? ??????
	DATA_IS_pix_ch_3	: out  std_logic_vector (bit_data_imx-1 downto 0);	-- ???????? ??????
	DATA_IS_pix_ch_4	: out  std_logic_vector (bit_data_imx-1 downto 0)	-- ???????? ??????
	);
end component;

signal DATA_IS_pix_ch_1		: std_logic_vector (bit_data_imx-1 downto 0);
signal DATA_IS_pix_ch_2		: std_logic_vector (bit_data_imx-1 downto 0);
signal DATA_IS_pix_ch_3		: std_logic_vector (bit_data_imx-1 downto 0);
signal DATA_IS_pix_ch_4		: std_logic_vector (bit_data_imx-1 downto 0);
----------------------------------------------------------------------


----------------------------------------------------------------------
-- ?????? ????????? ???????????? ?? ????????????? ????? ?????????????
----------------------------------------------------------------------
component IS_SIM_serial_DDR is
generic  (bit_data	: integer);
port (
		--??????? ???????--	
	CLK_fast				: in std_logic;  												-- ???????? 
	main_reset			: in std_logic;  												-- main_reset
	main_enable			: in std_logic;  												-- main_enable
	DATA_IMX_OUT		: in std_logic_vector (bit_data_imx-1 downto 0);	-- ??????? ??????
		--???????? ???????--	
	IMX_DDR_VIDEO		: out std_logic												-- ???????? ??????
		);
end component;
------------------------------------------------------------------------------------

begin
----------------------------------------------------------------------
-- ?????? PLL ??? ??????????? ?????? ?? ?????????????
-- ----------------------------------------------------------------------
-- PLL_POWERDOWN_N	<=	'1';
-- PLL_SIM_IS_q0: PLL_SIM_IS                   
-- port map (
-- 	-- Inputs
-- 	POWERDOWN	=> PLL_POWERDOWN_N,
-- 	CLKA			=> CLK,				--74.25 ???
-- 	-- Outputs 
-- 	GLA			=> CLK_IS_pix,		--137.5 ???
-- 	LOCK			=> locked_pll_0
-- );	
-- PLL_SIM_IS_q1: PLL_SIM_IS_1                   
-- port map (
-- 	-- Inputs
-- 	POWERDOWN	=> PLL_POWERDOWN_N,
-- 	CLKA			=> CLK,				--74.25 ???
-- 	-- Outputs 
-- 	GLA			=> CLK_IS_DDR_0, 	--206.25 ???	// ? ?????? LVDS 4 ch 12 bit
-- 	GLB			=> CLK_IS_DDR_1, 	--206.25 ???	// 180 phase shift
-- 	GLC			=> CLK_IS_DDR_2, 	--206.25 ???	// 90 phase shift
-- 	LOCK			=> locked_pll_1
-- );	


-- XVS_Imx_Sim <=	CLK_IS_pix;		
-- XHS_Imx_Sim	<=	CLK_IS_DDR_0;			
-- DATA_IS_PAR	<=	CLK_IS_DDR_1;			
-- DATA_IS_LVDS_ch_n<=	CLK_IS_DDR_2;		
-- DATA_IS_CSI	<=	locked_pll_1;			
-- CLK_DDR		<=	CLK_IS_pix;			
XVS_Imx_Sim <=	CLK;		
XHS_Imx_Sim	<=	CLK;			
-- DATA_IS_PAR	<=	CLK;			
-- DATA_IS_LVDS_ch_n<=	CLK;		
DATA_IS_CSI	<=	CLK;			
CLK_DDR		<=	CLK;			



-- ----------------------------------------------------------------------
-- -- ???????? reset ??? ??????????? ?????? 
-- ----------------------------------------------------------------------
-- process (CLK)
-- begin
-- if  rising_edge(CLK) then
-- 	locked_pll_q(0) <= locked_pll_0 or locked_pll_1;
-- 	for i in 0 to 30 loop
-- 		locked_pll_q(i+1) <= locked_pll_q(i);
-- 	end loop;
-- 	main_reset	<=	not 	locked_pll_q(31);
-- 	main_enable	<=	locked_pll_q(31);
-- end if;
-- end process;

-- ----------------------------------------------------------------------
-- -- ?????? ????????? ???????????? ?? ????????????? ? ???????????? ????
-- ----------------------------------------------------------------------
-- IS_SIM_Paralell_q: IS_SIM_Paralell    
-- generic map (
-- 	-- EKD_2200_1250p50.PixPerLine,
-- 	-- EKD_2200_1250p50.HsyncShift,
-- 	-- EKD_2200_1250p50.ActivePixPerLine,
-- 	-- EKD_2200_1250p50.HsyncWidth,
-- 	-- EKD_2200_1250p50.LinePerFrame,
-- 	-- EKD_2200_1250p50.VsyncShift,
-- 	-- EKD_2200_1250p50.ActiveLine,
-- 	-- EKD_2200_1250p50.VsyncWidth

-- 	EKD_ADV7343_1080p25.PixPerLine,
-- 	EKD_ADV7343_1080p25.HsyncShift,
-- 	EKD_ADV7343_1080p25.ActivePixPerLine,
-- 	EKD_ADV7343_1080p25.HsyncWidth,
-- 	EKD_ADV7343_1080p25.LinePerFrame,
-- 	EKD_ADV7343_1080p25.VsyncShift,
-- 	EKD_ADV7343_1080p25.ActiveLine,
-- 	EKD_ADV7343_1080p25.VsyncWidth


-- 	)
-- port map (
-- 				------??????? ???????-----------
-- 	CLK					=>	CLK_IS_pix,			
-- 	main_reset			=>	main_reset ,
-- 	main_enable			=>	main_enable  ,		
-- 	mode_generator		=>	mode_generator,
-- 				------???????? ???????-----------
-- 	DATA_IS_pix_ch_1	=> DATA_IS_pix_ch_1,
-- 	DATA_IS_pix_ch_2	=> DATA_IS_pix_ch_2,
-- 	DATA_IS_pix_ch_3	=> DATA_IS_pix_ch_3,
-- 	DATA_IS_pix_ch_4	=> DATA_IS_pix_ch_4
-- 	);	
-- ----------------------------------------------------------------------
-- -- ?????? ????????? ???????????? ?? ????????????? ????? ?????????????
-- -- ?????? ????? ???????? ?????????????? ??????????
-- ----------------------------------------------------------------------
-- IS_SIM_serial_DDR_q1: IS_SIM_serial_DDR                   
-- generic map (bit_data_imx) 
-- port map (
-- 				------??????? ???????-----------
-- 	CLK_fast				=>	CLK_IS_DDR_0,			
-- 	main_reset			=>	main_reset ,
-- 	main_enable			=>	main_enable  ,		
-- 	DATA_IMX_OUT		=>	DATA_IS_pix_ch_1,
-- 				------???????? ???????-----------
-- 	IMX_DDR_VIDEO		=>	DATA_IS_LVDS_ch_n(0)
-- 	);	
-- IS_SIM_serial_DDR_q2: IS_SIM_serial_DDR                   
-- generic map (bit_data_imx) 
-- port map (
-- 				------??????? ???????-----------
-- 	CLK_fast				=>	CLK_IS_DDR_0,			
-- 	main_reset			=>	main_reset ,
-- 	main_enable			=>	main_enable  ,		
-- 	DATA_IMX_OUT		=>	DATA_IS_pix_ch_2,
-- 				------???????? ???????-----------
-- 	IMX_DDR_VIDEO		=>	DATA_IS_LVDS_ch_n(1)
-- 	);	
-- IS_SIM_serial_DDR_q3: IS_SIM_serial_DDR                   
-- generic map (bit_data_imx) 
-- port map (
-- 				------??????? ???????-----------
-- 	CLK_fast				=>	CLK_IS_DDR_0,			
-- 	main_reset			=>	main_reset ,
-- 	main_enable			=>	main_enable  ,		
-- 	DATA_IMX_OUT		=>	DATA_IS_pix_ch_3,
-- 				------???????? ???????-----------
-- 	IMX_DDR_VIDEO		=>	DATA_IS_LVDS_ch_n(2)
-- 	);	
-- IS_SIM_serial_DDR_q4: IS_SIM_serial_DDR                   
-- generic map (bit_data_imx) 
-- port map (
-- 				------??????? ???????-----------
-- 	CLK_fast				=>	CLK_IS_DDR_0,			
-- 	main_reset			=>	main_reset ,
-- 	main_enable			=>	main_enable  ,		
-- 	DATA_IMX_OUT		=>	DATA_IS_pix_ch_4,
-- 				------???????? ???????-----------
-- 	IMX_DDR_VIDEO		=>	DATA_IS_LVDS_ch_n(3)
-- 	);	

-- CLK_DDR	<=	CLK_IS_DDR_2;

end ;
